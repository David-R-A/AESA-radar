library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.devkit_lib.all;

package params_pkg is
	-- DBF Params
	constant DBF_PARAMS : complex_int_matrix(0 to nA-1, 0 to nB-1) := (
		0 => (
			0 => (r => "00000011000001011111", i => "11111101011000011000"),
			1 => (r => "11111100011110011010", i => "11111110000111000000"),
			2 => (r => "11111101010001110101", i => "00000010111011100111"),
			3 => (r => "11111111101010101010", i => "00000011111111000111"),
			4 => (r => "11111111101010101010", i => "00000011111111000111"),
			5 => (r => "11111101010001110101", i => "00000010111011100111"),
			6 => (r => "11111100011110011010", i => "11111110000111000000"),
			7 => (r => "00000011000001011111", i => "11111101011000011000")
		),
		1 => (
			0 => (r => "11111101110101111011", i => "00000100101000010111"),
			1 => (r => "00000100111010101010", i => "00000001011000110100"),
			2 => (r => "00000011001010111010", i => "11111011111111101000"),
			3 => (r => "00000000011000011001", i => "11111010111001111101"),
			4 => (r => "00000000011000011001", i => "11111010111001111101"),
			5 => (r => "00000011001010111010", i => "11111011111111101000"),
			6 => (r => "00000100111010101010", i => "00000001011000110100"),
			7 => (r => "11111101110101111011", i => "00000100101000010111")
		),
		2 => (
			0 => (r => "00000000000110110011", i => "11111000111101111111"),
			1 => (r => "11111000111110101100", i => "11111111100101111100"),
			2 => (r => "11111100000101010100", i => "00000101110101110011"),
			3 => (r => "11111111100010011000", i => "00000111000001000110"),
			4 => (r => "11111111100010011000", i => "00000111000001000110"),
			5 => (r => "11111100000101010100", i => "00000101110101110011"),
			6 => (r => "11111000111110101100", i => "11111111100101111100"),
			7 => (r => "00000000000110110011", i => "11111000111101111111")
		),
		3 => (
			0 => (r => "00000011101011110100", i => "00001000100100110111"),
			1 => (r => "00001001001101110101", i => "11111110100001010011"),
			2 => (r => "00000100100100101010", i => "11110111110111001110"),
			3 => (r => "00000000100010000110", i => "11110110101011100110"),
			4 => (r => "00000000100010000110", i => "11110110101011100110"),
			5 => (r => "00000100100100101010", i => "11110111110111001110"),
			6 => (r => "00001001001101110101", i => "11111110100001010011"),
			7 => (r => "00000011101011110100", i => "00001000100100110111")
		),
		4 => (
			0 => (r => "11110111011101011100", i => "11111000001000110011"),
			1 => (r => "11110101001101000101", i => "00000100010001000101"),
			2 => (r => "11111011001000001000", i => "00001010100010010011"),
			3 => (r => "11111111011100001000", i => "00001011100110000100"),
			4 => (r => "11111111011100001000", i => "00001011100110000100"),
			5 => (r => "11111011001000001000", i => "00001010100010010011"),
			6 => (r => "11110101001101000101", i => "00000100010001000101"),
			7 => (r => "11110111011101011100", i => "11111000001000110011")
		),
		5 => (
			0 => (r => "00001100110111000011", i => "00000100010011101100"),
			1 => (r => "00001011001111100010", i => "11111000011010100010"),
			2 => (r => "00000100101101010000", i => "11110011010001111110"),
			3 => (r => "00000000100010010011", i => "11110010011100101100"),
			4 => (r => "00000000100010010011", i => "11110010011100101100"),
			5 => (r => "00000100101101010000", i => "11110011010001111110"),
			6 => (r => "00001011001111100010", i => "11111000011010100010"),
			7 => (r => "00001100110111000011", i => "00000100010011101100")
		),
		6 => (
			0 => (r => "11110001000100111011", i => "00000001011101100101"),
			1 => (r => "11110101101010110101", i => "00001010110111100010"),
			2 => (r => "11111011111010110010", i => "00001110011011011010"),
			3 => (r => "11111111100010100000", i => "00001110111111001100"),
			4 => (r => "11111111100010100000", i => "00001110111111001100"),
			5 => (r => "11111011111010110010", i => "00001110011011011010"),
			6 => (r => "11110101101010110101", i => "00001010110111100010"),
			7 => (r => "11110001000100111011", i => "00000001011101100101")
		),
		7 => (
			0 => (r => "00001101101011110010", i => "11111000001100001111"),
			1 => (r => "00001000001000111101", i => "11110010100000101010"),
			2 => (r => "00000011000101010010", i => "11110000100011001001"),
			3 => (r => "00000000010110001001", i => "11110000001111111010"),
			4 => (r => "00000000010110001001", i => "11110000001111111010"),
			5 => (r => "00000011000101010010", i => "11110000100011001001"),
			6 => (r => "00001000001000111101", i => "11110010100000101010"),
			7 => (r => "00001101101011110010", i => "11111000001100001111")
		),
		8 => (
			0 => (r => "11110110101100110110", i => "00001100101101111110"),
			1 => (r => "11111010111101010100", i => "00001110111011010100"),
			2 => (r => "11111110001001001001", i => "00001111101001010100"),
			3 => (r => "11111111110010101110", i => "00001111110000010000"),
			4 => (r => "11111111110010101110", i => "00001111110000010000"),
			5 => (r => "11111110001001001001", i => "00001111101001010100"),
			6 => (r => "11111010111101010100", i => "00001110111011010100"),
			7 => (r => "11110110101100110110", i => "00001100101101111110")
		),
		9 => (
			0 => (r => "00000011001000011110", i => "11110001010101100010"),
			1 => (r => "00000001101000000000", i => "11110001000110000001"),
			2 => (r => "00000000100101110010", i => "11110001000001000111"),
			3 => (r => "00000000000100001101", i => "11110001000000010111"),
			4 => (r => "00000000000100001101", i => "11110001000000010111"),
			5 => (r => "00000000100101110010", i => "11110001000001000111"),
			6 => (r => "00000001101000000000", i => "11110001000110000001"),
			7 => (r => "00000011001000011110", i => "11110001010101100010")
		),
		10 => (
			0 => (r => "00000010110101010101", i => "00001101010000110110"),
			1 => (r => "00000001011110000100", i => "00001101011110111000"),
			2 => (r => "00000000100010001011", i => "00001101100011010100"),
			3 => (r => "00000000000011110100", i => "00001101100011111111"),
			4 => (r => "00000000000011110100", i => "00001101100011111111"),
			5 => (r => "00000000100010001011", i => "00001101100011010100"),
			6 => (r => "00000001011110000100", i => "00001101011110111000"),
			7 => (r => "00000010110101010101", i => "00001101010000110110")
		),
		11 => (
			0 => (r => "11111001001001100000", i => "11110110101000010010"),
			1 => (r => "11111100010010010000", i => "11110101000000001001"),
			2 => (r => "11111110101000011011", i => "11110100011110010000"),
			3 => (r => "11111111110110001101", i => "11110100011001001001"),
			4 => (r => "11111111110110001101", i => "11110100011001001001"),
			5 => (r => "11111110101000011011", i => "11110100011110010000"),
			6 => (r => "11111100010010010000", i => "11110101000000001001"),
			7 => (r => "11111001001001100000", i => "11110110101000010010")
		),
		12 => (
			0 => (r => "00001000000110110110", i => "00000100101000000101"),
			1 => (r => "00000100110100101000", i => "00000111111111011110"),
			2 => (r => "00000001110100111000", i => "00001001001001110101"),
			3 => (r => "00000000001101000111", i => "00001001010101001111"),
			4 => (r => "00000000001101000111", i => "00001001010101001111"),
			5 => (r => "00000001110100111000", i => "00001001001001110101"),
			6 => (r => "00000100110100101000", i => "00000111111111011110"),
			7 => (r => "00001000000110110110", i => "00000100101000000101")
		),
		13 => (
			0 => (r => "11111001000000000101", i => "11111111010100000111"),
			1 => (r => "11111011001001111010", i => "11111010111001110011"),
			2 => (r => "11111110000101011111", i => "11111001001110111100"),
			3 => (r => "11111111110010001010", i => "11111000111110001001"),
			4 => (r => "11111111110010001010", i => "11111000111110001001"),
			5 => (r => "11111110000101011111", i => "11111001001110111100"),
			6 => (r => "11111011001001111010", i => "11111010111001110011"),
			7 => (r => "11111001000000000101", i => "11111111010100000111")
		),
		14 => (
			0 => (r => "00000100110110000001", i => "11111110011000001010"),
			1 => (r => "00000100001111000010", i => "00000010110110110111"),
			2 => (r => "00000001110001011110", i => "00000100110010101000"),
			3 => (r => "00000000001100111011", i => "00000101000110101101"),
			4 => (r => "00000000001100111011", i => "00000101000110101101"),
			5 => (r => "00000001110001011110", i => "00000100110010101000"),
			6 => (r => "00000100001111000010", i => "00000010110110110111"),
			7 => (r => "00000100110110000001", i => "11111110011000001010")
		),
		15 => (
			0 => (r => "11111101000011101011", i => "00000010101101011001"),
			1 => (r => "11111100010001111011", i => "11111110100001111010"),
			2 => (r => "11111110010100100010", i => "11111100010111101010"),
			3 => (r => "11111111110011101001", i => "11111100000000010011"),
			4 => (r => "11111111110011101001", i => "11111100000000010011"),
			5 => (r => "11111110010100100010", i => "11111100010111101010"),
			6 => (r => "11111100010001111011", i => "11111110100001111010"),
			7 => (r => "11111101000011101011", i => "00000010101101011001")
		)
	);

	-- PC Params
	constant PC_PARAMS : complex_in_vector(0 to PC_TAPS-1) := (
		0 => (r => "0000000000000000", i => "0000000000000000"),
		1 => (r => "0000110011001101", i => "0000110011001101"),
		2 => (r => "0001100110011010", i => "0001100110011010"),
		3 => (r => "0000110011001101", i => "0000110011001101"),
		4 => (r => "0000000000000000", i => "0000000000000000")
	);
end package params_pkg;